localparam  Z3_IDLE  = 2'd0,
            Z3_START = 2'd1,
            Z3_DATA  = 2'd2,
            Z3_END   = 2'd3;